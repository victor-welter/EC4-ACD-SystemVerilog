/**
*Codigo teste de modulo Aula2
*
*Autor: Víctor Vinicius Welter
*
*Data: Agosto de 2022
*
*Especificacao:
*Modulo teste
*/

module exe_01 (
    input logic in1,
    input logic in2,
    input logic in3,

    output logic out1,
    output logic out2
    
);
    
endmodule