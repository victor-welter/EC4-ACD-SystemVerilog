package definitions;
    typedef logic [15:0] word_t;
    typedef logic [31:0] dword_t; 
endpackage